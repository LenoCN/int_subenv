`ifndef INT_INTERFACE1
`define INT_INTERFACE1

interface int_interface;

    logic [31:0] test_signal = 'hABCD_1234;

endinterface

`endif
