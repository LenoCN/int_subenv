// IO Die interrupt entries to be added to int_map_entries.svh
// Generated based on IOSUB中断源 worksheet and SCP M7 interrupt list

        entry = '{name:"io_die_intr_0_intr", index:0, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[0]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[62]", dest_index_scp:62, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_1_intr", index:1, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[1]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[63]", dest_index_scp:63, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_2_intr", index:2, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[2]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[64]", dest_index_scp:64, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_3_intr", index:3, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[3]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[65]", dest_index_scp:65, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_4_intr", index:4, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[4]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[66]", dest_index_scp:66, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_5_intr", index:5, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[5]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[67]", dest_index_scp:67, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_6_intr", index:6, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[6]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[68]", dest_index_scp:68, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_7_intr", index:7, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[7]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[69]", dest_index_scp:69, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_8_intr", index:8, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[8]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[70]", dest_index_scp:70, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_9_intr", index:9, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[9]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[71]", dest_index_scp:71, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_10_intr", index:10, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[10]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[72]", dest_index_scp:72, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_11_intr", index:11, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[11]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[73]", dest_index_scp:73, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_12_intr", index:12, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[12]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[74]", dest_index_scp:74, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_13_intr", index:13, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[13]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[75]", dest_index_scp:75, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_14_intr", index:14, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[14]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[76]", dest_index_scp:76, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_15_intr", index:15, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[15]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[77]", dest_index_scp:77, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_16_intr", index:16, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[16]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[78]", dest_index_scp:78, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_17_intr", index:17, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[17]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[79]", dest_index_scp:79, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_18_intr", index:18, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[18]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[80]", dest_index_scp:80, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_19_intr", index:19, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[19]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[81]", dest_index_scp:81, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_20_intr", index:20, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[20]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[82]", dest_index_scp:82, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_21_intr", index:21, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[21]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[83]", dest_index_scp:83, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_22_intr", index:22, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[22]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[84]", dest_index_scp:84, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_23_intr", index:23, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[23]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[85]", dest_index_scp:85, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_24_intr", index:24, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[24]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[86]", dest_index_scp:86, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_25_intr", index:25, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[25]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[87]", dest_index_scp:87, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_26_intr", index:26, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[26]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[88]", dest_index_scp:88, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_27_intr", index:27, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[27]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[89]", dest_index_scp:89, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_28_intr", index:28, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[28]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[90]", dest_index_scp:90, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_29_intr", index:29, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[29]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[91]", dest_index_scp:91, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_30_intr", index:30, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[30]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[92]", dest_index_scp:92, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"io_die_intr_31_intr", index:31, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[31]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[93]", dest_index_scp:93, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);

// Total 32 IO Die interrupt entries generated
