`ifndef INT_ROUTING_MODEL_SV
`define INT_ROUTING_MODEL_SV

`include "int_def.sv"

// This class serves as the prediction model for interrupt routing.
// It is populated with data parsed from '中断向量表-iosub-V0.5.csv'.
class int_routing_model;
    
    // The main data structure holding all interrupt information.
    static interrupt_info_s interrupt_map[];

    // `build` function to populate the interrupt map.
    // NOTE: RTL paths are placeholders and need to be updated based on the final RTL hierarchy from int_harness.sv
    static function void build();
        interrupt_info_s entry;
        interrupt_group_e current_group;

        if (interrupt_map.size() > 0) return; // a simple guard to prevent multiple builds

        // --- Start of IOSUB interrupts ---
        current_group = IOSUB;
        entry = '{name:"iosub_slv_err_intr", index:0, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 0), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 0), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_buffer_ovf_intr", index:1, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 1), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 1), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_timeout_intr", index:2, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 2), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 2), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_qspi_intr", index:3, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 3), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 3), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 3), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_spi_intr", index:4, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 4), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 4), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 4), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_i2c0_intr", index:5, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 5), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 5), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_i2c1_intr", index:6, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 6), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 6), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_i2c2_intr", index:7, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 7), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 7), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pmbus0_intr", index:8, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 8), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:1, rtl_path_other_die:$sformatf("top_tb.int_harness.u_dut.other_die_bus[%0d]", 8)}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pmbus1_intr", index:9, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 9), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_uart0_intr", index:10, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 10), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 10), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_uart1_intr", index:11, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 11), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 11), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 11), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_uart2_intr", index:12, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 12), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 12), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 12), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_uart3_intr", index:13, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 13), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 13), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 13), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_uart4_intr", index:14, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 14), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 14), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 14), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dimm_i3c0_intr", index:15, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 15), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 15), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dimm_i3c1_intr", index:16, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 16), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 16), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dimm_i3c2_intr", index:17, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 17), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 17), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_sideband_i3c0_intr", index:18, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 18), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 18), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_gpio0_intr", index:19, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 19), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 19), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_gpio1_intr", index:20, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 20), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 20), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_gpio2_intr", index:21, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 21), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 21), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii0_q0_intr", index:22, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 22), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 22), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii0_q1_intr", index:23, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 23), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 23), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii0_q2_intr", index:24, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 24), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 24), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii0_q3_intr", index:25, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 25), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 25), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii1_q0_intr", index:26, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 26), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 26), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii1_q1_intr", index:27, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 27), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 27), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii1_q2_intr", index:28, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 28), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 28), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_rgmii1_q3_intr", index:29, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 29), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 29), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pvt_intr", index:30, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 30), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 30), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:1, rtl_path_other_die:$sformatf("top_tb.int_harness.u_dut.other_die_bus[%0d]", 30)}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dfx_lte_intr", index:31, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 31), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 31), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dw_axi_dlock_intr", index:32, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 32), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 32), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_mem_ist_intr", index:33, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 33), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_comreg_intr", index:34, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 34), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 34), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 34), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch0_intr", index:35, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 35), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 35), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 35), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch1_intr", index:36, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 36), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 36), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 36), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch2_intr", index:37, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 37), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 37), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 37), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch3_intr", index:38, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 38), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 38), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 38), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch4_intr", index:39, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 39), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 39), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 39), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch5_intr", index:40, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 40), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 40), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 40), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch6_intr", index:41, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 41), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 41), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 41), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch7_intr", index:42, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 42), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 42), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 42), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch8_intr", index:43, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 43), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 43), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 43), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch9_intr", index:44, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 44), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 44), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 44), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch10_intr", index:45, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 45), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 45), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 45), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch11_intr", index:46, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 46), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 46), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 46), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch12_intr", index:47, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 47), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 47), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 47), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch13_intr", index:48, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 48), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 48), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 48), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch14_intr", index:49, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 49), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 49), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 49), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_dma_ch15_intr", index:50, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 50), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 50), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 50), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_0_intr", index:51, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 51), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 51), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 51), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 51), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 51), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_1_intr", index:52, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 52), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 52), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 52), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 52), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 52), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_2_intr", index:53, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 53), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 53), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 53), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 53), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 53), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_3_intr", index:54, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 54), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 54), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 54), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 54), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 54), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_4_intr", index:55, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 55), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 55), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 55), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 55), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 55), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_5_intr", index:56, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 56), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 56), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 56), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 56), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 56), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_6_intr", index:57, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 57), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 57), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 57), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 57), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 57), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_7_intr", index:58, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 58), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 58), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 58), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 58), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 58), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_8_intr", index:59, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 59), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 59), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 59), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 59), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 59), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_9_intr", index:60, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 60), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 60), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 60), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 60), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 60), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_10_intr", index:61, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 61), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 61), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 61), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 61), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 61), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_11_intr", index:62, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 62), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 62), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 62), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 62), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 62), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_12_intr", index:63, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 63), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 63), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 63), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 63), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 63), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_13_intr", index:64, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 64), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 64), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 64), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 64), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 64), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_14_intr", index:65, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 65), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 65), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 65), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 65), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 65), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pad_in_15_intr", index:66, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 66), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 66), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 66), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 66), to_imu:1, rtl_path_imu:$sformatf("top_tb.int_harness.u_dut.imu_bus[%0d]", 66), to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_watchdog_io_intr", index:67, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 67), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 67), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 67), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 67), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pll_lock_intr", index:68, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 68), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_pll_unlock_intr", index:69, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 69), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_ras_cri_intr", index:70, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 70), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 70), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 70), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 70), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_ras_eri_intr", index:71, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 71), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 71), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 71), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 71), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_ras_fhi_intr", index:72, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 72), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 72), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 72), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 72), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_strap_load_fail_intr", index:73, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 73), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:1, rtl_path_io:$sformatf("top_tb.int_harness.u_dut.io_bus[%0d]", 73), to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_abnormal_0_intr", index:74, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 74), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 74), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 74), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 74), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_abnormal_1_intr", index:75, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 75), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 75), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 75), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 75), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"iosub_normal_intr", index:76, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 76), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 76), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 76), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"pvt_temp_alarm_intr", index:77, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 77), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:1, rtl_path_io:$sformatf("top_tb.int_harness.u_dut.io_bus[%0d]", 77), to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"merge_pll_intr_lock", index:78, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 78), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 78), to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"merge_pll_intr_unlock", index:79, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 79), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 79), to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"merge_pll_intr_frechangedone", index:80, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 80), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 80), to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"merge_pll_intr_frechange_tot_done", index:81, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 81), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 81), to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"merge_pll_intr_intdocfrac_err", index:82, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.iosub_interrupts[%0d]", 82), to_ap:0, rtl_path_ap:"", to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 82), to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);

        // --- Start of USB interrupts ---
        current_group = USB;
        entry = '{name:"usb0_ctrl_xhci_intr", index:0, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 0), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 0), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb0_ctrl_otg_intr", index:1, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 1), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 1), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb0_ctrl_dev_intr", index:2, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 2), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 2), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb0_ctrl_sys_intr", index:3, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 3), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 3), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb0_phy3_intr", index:4, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 4), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 4), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_ctrl_xhci_intr", index:5, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 5), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 5), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_ctrl_otg_intr", index:6, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 6), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 6), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_ctrl_dev_intr", index:7, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 7), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 7), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_ctrl_sys_intr", index:8, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 8), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 8), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_phy3_intr", index:9, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 9), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 9), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb0_apb1ton_intr", index:10, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 10), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb1_apb1ton_intr", index:11, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 11), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"usb_top_apb1ton_intr", index:12, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.usb_interrupts[%0d]", 12), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);

        // --- Start of SMMU interrupts ---
        current_group = SMMU;
        entry = '{name:"intr_tcu_ups_event_q_irpt_s", index:0, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 0), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 0), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_cmd_sync_irpt_s", index:1, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 1), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 1), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_global_irpt_s", index:2, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 2), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 2), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_gpf_far", index:3, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 3), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 3), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_gpt_cfg_far", index:4, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 4), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 4), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_event_q_irpt_ns", index:5, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 5), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 5), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_cmd_sync_irpt_ns", index:6, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 6), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 6), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_global_irpt_ns", index:7, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 7), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 7), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_pmu_irpt", index:8, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 8), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 8), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tcu_ups_pri_q_irpt_ns", index:9, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 9), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 9), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tbu0_ups_pmu_irpt", index:10, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 10), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 10), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"intr_tbu0_ups_crit_err", index:11, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 11), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 11), to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_abnormal_intr", index:12, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 12), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 12), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 12), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 12), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_normal_intr_ns", index:13, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 13), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 13), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 13), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 13), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_normal_intr_s", index:14, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 14), to_ap:1, rtl_path_ap:$sformatf("top_tb.int_harness.u_dut.ap_bus[%0d]", 14), to_scp:1, rtl_path_scp:$sformatf("top_tb.int_harness.u_dut.scp_bus[%0d]", 14), to_mcp:1, rtl_path_mcp:$sformatf("top_tb.int_harness.u_dut.mcp_bus[%0d]", 14), to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_cri_intr", index:15, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 15), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_eri_intr", index:16, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 16), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);
        entry = '{name:"smmu_fhi_intr", index:17, group:current_group, rtl_path_src:$sformatf("top_tb.int_harness.u_dut.smmu_interrupts[%0d]", 17), to_ap:0, rtl_path_ap:"", to_scp:0, rtl_path_scp:"", to_mcp:0, rtl_path_mcp:"", to_imu:0, rtl_path_imu:"", to_io:0, rtl_path_io:"", to_other_die:0, rtl_path_other_die:""}; interrupt_map.push_back(entry);

        // --- Add more groups as needed based on CSV ---
        // TODO: Populate other interrupt groups (SCP, MCP, IODAP, etc.) in a similar fashion.
    endfunction

endclass

`endif // INT_ROUTING_MODEL_SV
