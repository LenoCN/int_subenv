// Missing interrupt entries to be added to int_map_entries.svh
// Generated based on IOSUB中断源 worksheet and SCP/MCP M7 interrupt lists

        entry = '{name:"ap2scp_mhu_receive_intr_0", index:32, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[32]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[32]", dest_index_scp:32, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"ap2scp_mhu_receive_intr_1", index:33, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[33]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[33]", dest_index_scp:33, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"ap2scp_mhu_receive_intr_2", index:34, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[34]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[34]", dest_index_scp:34, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"ap2scp_mhu_receive_intr_3", index:35, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[35]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[35]", dest_index_scp:35, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d0_iosub_pmbus0_intr", index:97, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[97]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[52]", dest_index_scp:52, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d0_iosub_pvt_intr", index:98, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[98]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[53]", dest_index_scp:53, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d0_n2_wakeup_intr", index:95, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[95]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[50]", dest_index_scp:50, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d0_n2_ws1_intr", index:96, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[96]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[51]", dest_index_scp:51, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d1_iosub_pmbus0_intr", index:101, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[101]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[56]", dest_index_scp:56, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d1_iosub_pvt_intr", index:102, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[102]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[57]", dest_index_scp:57, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d1_n2_wakeup_intr", index:99, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[99]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[54]", dest_index_scp:54, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d1_n2_ws1_intr", index:100, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[100]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[55]", dest_index_scp:55, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d2_iosub_pmbus0_intr", index:105, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[105]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[60]", dest_index_scp:60, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d2_iosub_pvt_intr", index:106, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[106]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[61]", dest_index_scp:61, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d2_n2_wakeup_intr", index:103, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[103]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[58]", dest_index_scp:58, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_d2_n2_ws1_intr", index:104, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[104]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[59]", dest_index_scp:59, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_mcp2scp_mhu_receive_intr_0", index:69, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[69]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[47]", dest_index_scp:47, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_mcp2scp_mhu_receive_intr_1", index:70, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[70]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[48]", dest_index_scp:48, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_mcp2scp_mhu_receive_intr_2", index:71, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[71]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[49]", dest_index_scp:49, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2mcp_mhu_send_intr_0", index:51, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[51]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[41]", dest_index_scp:41, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2mcp_mhu_send_intr_1", index:52, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[52]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[42]", dest_index_scp:42, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2mcp_mhu_send_intr_2", index:53, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[53]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[43]", dest_index_scp:43, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_receive_intr_0", index:60, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[60]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[44]", dest_index_scp:44, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_receive_intr_1", index:61, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[61]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[45]", dest_index_scp:45, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_receive_intr_2", index:62, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[62]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[46]", dest_index_scp:46, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_send_intr_0", index:48, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[48]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[38]", dest_index_scp:38, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_send_intr_1", index:49, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[49]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[39]", dest_index_scp:39, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"d2d_scp2scp_mhu_send_intr_2", index:50, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[50]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[40]", dest_index_scp:40, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);

        entry = '{name:"mcp2io_wdt_ws1_intr", index:19, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[19]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp2scp_mhu_receive_intr", index:47, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[47]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[37]", dest_index_scp:37, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_acl_intr", index:13, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[13]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[10]", dest_index_mcp:10, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_cpu_bus_fault_intr", index:12, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[12]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[9]", dest_index_mcp:9, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_cpu_cti_irq[0]", index:14, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[14]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[11]", dest_index_mcp:11, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_cpu_cti_irq[1]", index:15, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[15]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[12]", dest_index_mcp:12, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_gpio_intr", index:10, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[10]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[7]", dest_index_mcp:7, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_i2c_intr", index:11, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[11]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[8]", dest_index_mcp:8, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_smbus_intr", index:9, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[9]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[6]", dest_index_mcp:6, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_sram_bus_fault_intr", index:20, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[20]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[13]", dest_index_mcp:13, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_timer64_0_intr", index:4, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[4]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[1]", dest_index_mcp:1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_timer64_1_intr", index:5, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[5]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[2]", dest_index_mcp:2, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_timer64_2_intr", index:6, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[6]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[3]", dest_index_mcp:3, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_timer64_3_intr", index:7, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[7]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[4]", dest_index_mcp:4, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"mcp_uart_intr", index:8, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[8]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:1, rtl_path_mcp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_mcp_top.u_cortexm7_wrapper.cpu_irq[5]", dest_index_mcp:5, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2ap_mhu_send_intr_0", index:12, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[12]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[28]", dest_index_scp:28, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2ap_mhu_send_intr_1", index:13, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[13]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[29]", dest_index_scp:29, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2ap_mhu_send_intr_2", index:14, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[14]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[30]", dest_index_scp:30, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2ap_mhu_send_intr_3", index:15, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[15]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[31]", dest_index_scp:31, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2io_wdt_ws1_intr", index:93, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[93]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:0, rtl_path_scp:"", dest_index_scp:-1, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp2mcp_mhu_send_intr", index:44, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[44]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[36]", dest_index_scp:36, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_acl_intr", index:9, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[9]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[6]", dest_index_scp:6, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_cpu_bus_fault_intr", index:8, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[8]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[5]", dest_index_scp:5, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_cpu_cti_irq[0]", index:10, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[10]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[7]", dest_index_scp:7, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_cpu_cti_irq[1]", index:11, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[11]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[8]", dest_index_scp:8, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_dma_intr", index:78, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[78]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[15]", dest_index_scp:15, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_efuse_intr", index:79, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[79]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[16]", dest_index_scp:16, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_gpio_intr", index:84, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[84]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[25]", dest_index_scp:25, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_i2c_intr", index:85, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[85]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[26]", dest_index_scp:26, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_i3c_dma_0_intr", index:75, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[75]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[12]", dest_index_scp:12, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_i3c_dma_1_intr", index:76, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[76]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[13]", dest_index_scp:13, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_i3c_dma_2_intr", index:77, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[77]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[14]", dest_index_scp:14, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_qspi_intr", index:80, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[80]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[17]", dest_index_scp:17, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_smbus_intr", index:83, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[83]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[24]", dest_index_scp:24, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_spi_intr", index:81, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[81]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[18]", dest_index_scp:18, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_sram_bus_fault_intr", index:94, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[94]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[27]", dest_index_scp:27, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_timer64_0_intr", index:4, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[4]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[1]", dest_index_scp:1, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_timer64_1_intr", index:5, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[5]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[2]", dest_index_scp:2, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_timer64_2_intr", index:6, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[6]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[3]", dest_index_scp:3, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_timer64_3_intr", index:7, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[7]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[4]", dest_index_scp:4, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_ts_sync_0_intr", index:72, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[72]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[9]", dest_index_scp:9, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_ts_sync_1_intr", index:73, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[73]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[10]", dest_index_scp:10, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_ts_sync_2_intr", index:74, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[74]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[11]", dest_index_scp:11, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"scp_uart_intr", index:82, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[82]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[23]", dest_index_scp:23, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);
        entry = '{name:"slcm_fault_intr", index:110, group:IOSUB, trigger:LEVEL, polarity:ACTIVE_HIGH, rtl_path_src:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_iosub_int_sub.iosub_peri_intr[110]", pulse_width_ns:0, to_ap:0, rtl_path_ap:"", dest_index_ap:-1, to_scp:1, rtl_path_scp:"top_tb.multidie_top.DUT[0].u_str_top.u_iosub_top_wrap.u0_iosub_top_wrap_hd.u0_iosub_top_wrap_raw.u_scp_top_wrapper.u_scp_top.u_m7_wrapper.cpu_irq[94]", dest_index_scp:94, to_mcp:0, rtl_path_mcp:"", dest_index_mcp:-1, to_accel:0, rtl_path_accel:"", dest_index_accel:-1, to_io:0, rtl_path_io:"", dest_index_io:-1, to_other_die:0, rtl_path_other_die:"", dest_index_other_die:-1}; interrupt_map.push_back(entry);

// Total 89 missing interrupt entries generated
